*=========================================================
* VGID Sweep (PMOS, NBTI) -- FIXED, 2-column output
*=========================================================

.include "C:/Users/Lenovo/Documents/bsim4_analyzer_reliability/models/pmos130.sp"

.temp 85.0

M1 d g s b pmos130 W=1e-06 L=1.3e-07

Vd d 0 0
Vs s 0 1.2
Vb b 0 0
Vg g s 0

.dc Vg 0 -1.2 -0.005

.control
  set filetype=ascii
  run

  let VX = v(g)-v(s)
  let IY = abs(i(Vd))

  * ======== FIX ========
  * 出力を HCI と同じ 2 列構造に統一
  wrdata 130nm_nbti_pmos_12v_85c_t0s_vgid.dat VX IY
  * =====================

  quit
.endc

.end
