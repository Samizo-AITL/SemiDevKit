* ============================================================
*  VGID Template (NMOS / PMOS 共通)
*  BSIM4 DIM: Id–Vg Sweep
*  - Python 側から {{…}} が埋め込まれる前提
* ============================================================

{{MODEL_INCLUDE}}

* -------------------------
* Geometry / Temperature
* -------------------------
.param LCH = {{LCH}}
.param WCH = {{WCH}}
.temp {{TEMP}}

* -------------------------
* Terminal voltages
*   - NMOS : D = VDD, S = 0,   B = 0
*   - PMOS : D = 0,   S = VDD, B = VDD
*   （いずれも Python 側で {{D_VOLT}}, {{S_VOLT}}, {{B_VOLT}} を設定）
* -------------------------
Vd   d      0      {{D_VOLT}}
Vs   s      0      {{S_VOLT}}
Vb   b      0      {{B_VOLT}}

* Gate sweep source (gate vs source)
Vg   g      s      0

* MOS Device
*   - L/W はパラメータ LCH/WCH を使用
*   - {{MODEL_NAME}} は Python 側で L/W 専用モデル名に差し替え
M1  d  g  s  b  {{MODEL_NAME}}  L=LCH  W=WCH

.options post=2 nomod

* Vg を掃引（NMOS: 0→VDD, PMOS: 0→-VDD）
.dc Vg {{VG_START}} {{VG_STOP}} {{VG_STEP}}

.control
  set filetype=ascii
  run

  * -------------------------------------
  * VX = Vgs  (v(g) - v(s))
  * -------------------------------------
  let VX = v(g) - v(s)

  * -------------------------------------
  * Id (Drain→Source の向きを正方向に統一)
  *
  * NMOS:
  *   Source = 0V  → Id = -I(Vd)
  *
  * PMOS:
  *   Source = VDD → Id =  I(Vs)
  *
  * {{S_VOLT}} は Python 側で
  *   - NMOS: 0
  *   - PMOS: VDD
  * に置換される前提
  * -------------------------------------
  if ( {{S_VOLT}} == 0 )
    * NMOS
    let IY = -i(Vd)
  else
    * PMOS
    let IY =  i(Vs)
  end

  * -------------------------------------
  * CSV (ASCII) 出力
  *   1列目: VX (= Vgs)
  *   2列目: IY (= Id, Ds 向き正)
  * -------------------------------------
  wrdata {{CSV_PATH}}  VX  IY
  quit
.endc

.end
