*=========================================================
* VGID Sweep (NMOS)
*=========================================================

{{MODEL_INCLUDE}}

.temp {{TEMP}}

M1 d g s b {{MODEL_NAME}} W={{WCH}} L={{LCH}}

Vd d 0 {{D_VOLT}}
Vs s 0 {{S_VOLT}}
Vb b 0 {{B_VOLT}}
Vg g s 0

.dc Vg {{VG_START}} {{VG_STOP}} {{VG_STEP}}

.control
  set filetype=ascii
  run

  let VX = v(g)-v(s)
  let IY = abs(i(Vd))

  wrdata {{CSV_PATH}} VX IY
  quit
.endc

.end
