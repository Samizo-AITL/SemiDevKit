* =========================================================
*  BSIM4 Simplified Model — Education Use
* =========================================================

* ---------- NMOS ---------------
.model nmos130 nmos level=54
+ version = 4.8
+ toxref  = 2.3e-9
+ vth0    = 0.40
+ u0      = 0.013
+ vsat    = 1.5e6
+ rdsw    = 80
+ k1      = 0.50
+ k2      = -0.03
+ voff    = -0.05
+ nfactor = 1.3
