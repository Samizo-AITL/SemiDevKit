* =========================================================
*  BSIM4 Simplified Model — Education Use
* =========================================================

* ---------- PMOS ---------------
.model pmos130 pmos level=54
+ version = 4.8
+ toxref  = 2.3e-9
+ vth0    = -0.40
+ u0      = 0.006
+ vsat    = 1.0e6
+ rdsw    = 120
+ k1      = 0.50
+ k2      = -0.03
+ voff    = -0.05
+ nfactor = 1.3
