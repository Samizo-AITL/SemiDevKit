*=========================================================
* PMOS NBTI Stress + DC Extraction
*=========================================================

.include "{{MODEL_FILE}}"

.temp {{STRESS_TEMP}}

* PMOS device
M1 d g s b pmos130 L=0.13u W=1u

* Bias
Vd d 0 {{STRESS_VDS}}
Vg g 0 {{STRESS_VGS}}
Vs s 0 1.2
Vb b 0 0

* DC operating point
.op

.control
  set filetype=ascii
  run

  let IDLIN = abs(i(Vd))
  let IDSAT = abs(i(Vd))

  wrdata {{LOG_FILE}} 0 IDLIN IDSAT
  quit
.endc

.end
