* Paramus Physical Edition generated BSIM4 modelcard
.model paramus_nmos nmos level=54
+ vth0    = -0.14496568148224975
+ u0      = 0.009999999999999887
+ pclm    = 0.1000000000000002
+ eta0    = 0.05
+ dvt0    = 1.0
+ dvt1    = 0.5
+ nfactor = 1.5
+ toxm    = 2.2e-09
+ rdsw    = 200.0
+ vsat    = 100000.0
+ k1      = 0.6
+ k2      = -0.02
+ cgso    = 1e-10
+ cgdo    = 1e-10
