* ============================================================
*  VDID Template (NMOS / PMOS 共通)
*  BSIM4 DIM : Id–Vd (Drain sweep)
* ============================================================

{{MODEL_INCLUDE}}

.param LCH      = {{LCH}}
.param WCH      = {{WCH}}
.param VG_BIAS  = {{VG_BIAS}}

.temp {{TEMP}}

* -------------------------
* Terminal Bias
* -------------------------
* NMOS :
*   S = 0V
*   B = 0V
*   Drain sweep: 0 → +VDD
*
* PMOS :
*   S = VDD
*   B = VDD
*   Drain sweep: 0 → –VDD
* -------------------------

Vs     s      0     {{S_VOLT}}
Vb     b      0     {{B_VOLT}}

* Drain sweep source
VDSRC  d_int  s     {{VD_START}}

* Gate bias
Vg     g      s     {{VG_BIAS}}

* MOS Device
M1  d_int  g  s  b  {{MODEL_NAME}}  L=LCH  W=WCH

.options post=2 nomod
.dc VDSRC {{VD_START}} {{VD_STOP}} {{VD_STEP}}

.control
  set filetype=ascii
  run

  * ------------------------------------------------
  * Current / Voltage Definitions
  *
  *  Id (positive when flowing Drain → Source)
  *
  *  NMOS :
  *     Id = -I(VDSRC)
  *     Vds = V(d) - V(s)
  *
  *  PMOS :
  *     Id = +I(VDSRC)
  *     Vds = V(d) - V(s)   (負になるが Id と整合する）
  *
  *  → VX : Drain-Source Voltage (Vds)
  *  → IY : Drain current (positive = Drain→Source)
  * ------------------------------------------------

  if ( {{S_VOLT}} > 0 )
    * PMOS
    let VX =  v(d_int) - v(s)     ; Vd - Vs  (PMOSでは負になる)
    let IY =  i(VDSRC)            ; PMOS Id
  else
    * NMOS
    let VX =  v(d_int) - v(s)     ; Vd - Vs
    let IY = -i(VDSRC)            ; NMOS Id
  end

  * ------------------------------------------------
  * Save as ASCII CSV
  *   col1 : VX = Vds
  *   col2 : IY = Id (D → S 正方向)
  * ------------------------------------------------
  wrdata {{DAT_PATH}}  VX  IY

  quit
.endc

.end
